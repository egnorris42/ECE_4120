-- Elizabeth Norris
-- ECE 4120 - Project Phase 3
-- 04/29/2021
-- .vhd

library ieee, lcdf_vhdl;
use ieee.std_logic_1164.all; 
use IEEE.std_logic_arith.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity  is
	port();
	end ;
	
architecture _behavior of  is


end _behavior;